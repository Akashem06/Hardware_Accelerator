`define INSTRUCTION_WIDTH 32      // Instruction width (in bits)
`define DATA_WIDTH 32             // Data width (in bits)
`define ADDR_WIDTH 32             // Address width for memory
`define NUM_REGS 32               // Number of registers in the register file
`define NUM_MEMORY_CELLS 1024     // Number of cells in memory
