`include "global_defines.sv"

module pipeline_control 
import matrix_ops_pkg::*;
(
    input logic clk,
    input logic rst_n,

    // Instruction fetch stage interface
    input logic                          fetch_valid,
    input logic [`INSTRUCTION_WIDTH-1:0] fetch_pc,
    output logic                         fetch_stall,
    output logic                         fetch_flush,

    // Decode stage interface
    input logic                          decode_valid,
    input logic [`INSTRUCTION_WIDTH-1:0] decoded_instruction,
    input logic                          is_matrix_op,
    input matrix_op_t                    matrix_op_type,
    output logic                         decode_stall,
    output logic                         decode_flush,

    // Execute stage interface
    input  logic        execute_valid,
    input  logic [4:0]  execute_rd,      // Destination register of executing instruction
    input  logic        execute_wb_en,   // Writeback enable in Execute stage
    input  logic [4:0]  execute_rs1,     // Source register 1 (for hazard checking)
    input  logic [4:0]  execute_rs2,     // Source register 2
    input  logic        matrix_busy,     // Matrix unit busy signal (from accelerator)
    output logic        execute_stall,
    output logic        execute_flush,
    
    // Memory stage interface
    input  logic        mem_valid,
    input  logic [4:0]  mem_rd,
    input  logic        mem_wb_en,
    
    // Writeback stage interface
    input  logic        wb_valid,
    input  logic [4:0]  wb_rd,
    input  logic        wb_wb_en
);

//-------------------------------------------------------------------------
// Internal signals for hazard detection
//-------------------------------------------------------------------------
logic data_hazard;
logic structural_hazard;
logic control_hazard = 1'b0;
logic matrix_conflict;

endmodule
