`define WORD_SIZE 4               // Word size in bytes
`define INSTRUCTION_WIDTH 32      // Instruction width (in bits)
`define DATA_WIDTH 32             // Data width (in bits)
`define ADDR_WIDTH 32             // Address width for memory
`define NUM_REGS 16               // Number of registers in the register file
`define NUM_REGS_BIT_COUNT 4      // Number of bits used to store the number of regs
`define NUM_MEMORY_CELLS 1024     // Number of cells in memory
`define NUM_MATRIX_COLS_ROWS 16   // Number of matrix columns/rows supported
