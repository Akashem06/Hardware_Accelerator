`include "global_defines.sv"

/* verilator lint_off UNUSED */
module top (
    input logic clk,
    input logic rst,
    input logic rst_n
);

endmodule
