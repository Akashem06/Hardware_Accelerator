`ifndef RISCV_PKG_SV
`define RISCV_PKG_SV

package riscv_pkg;
    parameter XLEN = 32;    // RV32 ISA
    parameter ILEN = 32;    // Instruction length
endpackage

`endif